module simple(cOut,x1,x2);
input x1,x2;
output cOut;
wire x1,x2,cOut;
assign cOut = x1 & x2;
endmodule
